module top();
    
endmodule
