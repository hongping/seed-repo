module testbench();
    top dut();

    initial $display("hello world!\n");
endmodule
